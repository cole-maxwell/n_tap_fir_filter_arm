// arm_hps.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module arm_hps (
		input  wire        clk_clk,             //          clk.clk
		output wire [12:0] memory_mem_a,        //       memory.mem_a
		output wire [2:0]  memory_mem_ba,       //             .mem_ba
		output wire        memory_mem_ck,       //             .mem_ck
		output wire        memory_mem_ck_n,     //             .mem_ck_n
		output wire        memory_mem_cke,      //             .mem_cke
		output wire        memory_mem_cs_n,     //             .mem_cs_n
		output wire        memory_mem_ras_n,    //             .mem_ras_n
		output wire        memory_mem_cas_n,    //             .mem_cas_n
		output wire        memory_mem_we_n,     //             .mem_we_n
		output wire        memory_mem_reset_n,  //             .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,       //             .mem_dq
		inout  wire        memory_mem_dqs,      //             .mem_dqs
		inout  wire        memory_mem_dqs_n,    //             .mem_dqs_n
		output wire        memory_mem_odt,      //             .mem_odt
		output wire        memory_mem_dm,       //             .mem_dm
		input  wire        memory_oct_rzqin,    //             .oct_rzqin
		output wire [31:0] pio_display_export,  //  pio_display.export
		input  wire [15:0] pio_fpga2hps_export, // pio_fpga2hps.export
		output wire [15:0] pio_hps2fpga_export, // pio_hps2fpga.export
		input  wire [3:0]  pio_keys_export,     //     pio_keys.export
		output wire [9:0]  pio_led_export,      //      pio_led.export
		input  wire        reset_reset_n        //        reset.reset_n
	);

	wire   [1:0] cpu_h2f_axi_master_awburst;                   // cpu:h2f_AWBURST -> mm_interconnect_0:cpu_h2f_axi_master_awburst
	wire   [3:0] cpu_h2f_axi_master_arlen;                     // cpu:h2f_ARLEN -> mm_interconnect_0:cpu_h2f_axi_master_arlen
	wire   [3:0] cpu_h2f_axi_master_wstrb;                     // cpu:h2f_WSTRB -> mm_interconnect_0:cpu_h2f_axi_master_wstrb
	wire         cpu_h2f_axi_master_wready;                    // mm_interconnect_0:cpu_h2f_axi_master_wready -> cpu:h2f_WREADY
	wire  [11:0] cpu_h2f_axi_master_rid;                       // mm_interconnect_0:cpu_h2f_axi_master_rid -> cpu:h2f_RID
	wire         cpu_h2f_axi_master_rready;                    // cpu:h2f_RREADY -> mm_interconnect_0:cpu_h2f_axi_master_rready
	wire   [3:0] cpu_h2f_axi_master_awlen;                     // cpu:h2f_AWLEN -> mm_interconnect_0:cpu_h2f_axi_master_awlen
	wire  [11:0] cpu_h2f_axi_master_wid;                       // cpu:h2f_WID -> mm_interconnect_0:cpu_h2f_axi_master_wid
	wire   [3:0] cpu_h2f_axi_master_arcache;                   // cpu:h2f_ARCACHE -> mm_interconnect_0:cpu_h2f_axi_master_arcache
	wire         cpu_h2f_axi_master_wvalid;                    // cpu:h2f_WVALID -> mm_interconnect_0:cpu_h2f_axi_master_wvalid
	wire  [29:0] cpu_h2f_axi_master_araddr;                    // cpu:h2f_ARADDR -> mm_interconnect_0:cpu_h2f_axi_master_araddr
	wire   [2:0] cpu_h2f_axi_master_arprot;                    // cpu:h2f_ARPROT -> mm_interconnect_0:cpu_h2f_axi_master_arprot
	wire   [2:0] cpu_h2f_axi_master_awprot;                    // cpu:h2f_AWPROT -> mm_interconnect_0:cpu_h2f_axi_master_awprot
	wire  [31:0] cpu_h2f_axi_master_wdata;                     // cpu:h2f_WDATA -> mm_interconnect_0:cpu_h2f_axi_master_wdata
	wire         cpu_h2f_axi_master_arvalid;                   // cpu:h2f_ARVALID -> mm_interconnect_0:cpu_h2f_axi_master_arvalid
	wire   [3:0] cpu_h2f_axi_master_awcache;                   // cpu:h2f_AWCACHE -> mm_interconnect_0:cpu_h2f_axi_master_awcache
	wire  [11:0] cpu_h2f_axi_master_arid;                      // cpu:h2f_ARID -> mm_interconnect_0:cpu_h2f_axi_master_arid
	wire   [1:0] cpu_h2f_axi_master_arlock;                    // cpu:h2f_ARLOCK -> mm_interconnect_0:cpu_h2f_axi_master_arlock
	wire   [1:0] cpu_h2f_axi_master_awlock;                    // cpu:h2f_AWLOCK -> mm_interconnect_0:cpu_h2f_axi_master_awlock
	wire  [29:0] cpu_h2f_axi_master_awaddr;                    // cpu:h2f_AWADDR -> mm_interconnect_0:cpu_h2f_axi_master_awaddr
	wire   [1:0] cpu_h2f_axi_master_bresp;                     // mm_interconnect_0:cpu_h2f_axi_master_bresp -> cpu:h2f_BRESP
	wire         cpu_h2f_axi_master_arready;                   // mm_interconnect_0:cpu_h2f_axi_master_arready -> cpu:h2f_ARREADY
	wire  [31:0] cpu_h2f_axi_master_rdata;                     // mm_interconnect_0:cpu_h2f_axi_master_rdata -> cpu:h2f_RDATA
	wire         cpu_h2f_axi_master_awready;                   // mm_interconnect_0:cpu_h2f_axi_master_awready -> cpu:h2f_AWREADY
	wire   [1:0] cpu_h2f_axi_master_arburst;                   // cpu:h2f_ARBURST -> mm_interconnect_0:cpu_h2f_axi_master_arburst
	wire   [2:0] cpu_h2f_axi_master_arsize;                    // cpu:h2f_ARSIZE -> mm_interconnect_0:cpu_h2f_axi_master_arsize
	wire         cpu_h2f_axi_master_bready;                    // cpu:h2f_BREADY -> mm_interconnect_0:cpu_h2f_axi_master_bready
	wire         cpu_h2f_axi_master_rlast;                     // mm_interconnect_0:cpu_h2f_axi_master_rlast -> cpu:h2f_RLAST
	wire         cpu_h2f_axi_master_wlast;                     // cpu:h2f_WLAST -> mm_interconnect_0:cpu_h2f_axi_master_wlast
	wire   [1:0] cpu_h2f_axi_master_rresp;                     // mm_interconnect_0:cpu_h2f_axi_master_rresp -> cpu:h2f_RRESP
	wire  [11:0] cpu_h2f_axi_master_awid;                      // cpu:h2f_AWID -> mm_interconnect_0:cpu_h2f_axi_master_awid
	wire  [11:0] cpu_h2f_axi_master_bid;                       // mm_interconnect_0:cpu_h2f_axi_master_bid -> cpu:h2f_BID
	wire         cpu_h2f_axi_master_bvalid;                    // mm_interconnect_0:cpu_h2f_axi_master_bvalid -> cpu:h2f_BVALID
	wire   [2:0] cpu_h2f_axi_master_awsize;                    // cpu:h2f_AWSIZE -> mm_interconnect_0:cpu_h2f_axi_master_awsize
	wire         cpu_h2f_axi_master_awvalid;                   // cpu:h2f_AWVALID -> mm_interconnect_0:cpu_h2f_axi_master_awvalid
	wire         cpu_h2f_axi_master_rvalid;                    // mm_interconnect_0:cpu_h2f_axi_master_rvalid -> cpu:h2f_RVALID
	wire         mm_interconnect_0_ram_s1_chipselect;          // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;            // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;             // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;          // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;               // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;           // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;               // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire   [1:0] cpu_h2f_lw_axi_master_awburst;                // cpu:h2f_lw_AWBURST -> mm_interconnect_1:cpu_h2f_lw_axi_master_awburst
	wire   [3:0] cpu_h2f_lw_axi_master_arlen;                  // cpu:h2f_lw_ARLEN -> mm_interconnect_1:cpu_h2f_lw_axi_master_arlen
	wire   [3:0] cpu_h2f_lw_axi_master_wstrb;                  // cpu:h2f_lw_WSTRB -> mm_interconnect_1:cpu_h2f_lw_axi_master_wstrb
	wire         cpu_h2f_lw_axi_master_wready;                 // mm_interconnect_1:cpu_h2f_lw_axi_master_wready -> cpu:h2f_lw_WREADY
	wire  [11:0] cpu_h2f_lw_axi_master_rid;                    // mm_interconnect_1:cpu_h2f_lw_axi_master_rid -> cpu:h2f_lw_RID
	wire         cpu_h2f_lw_axi_master_rready;                 // cpu:h2f_lw_RREADY -> mm_interconnect_1:cpu_h2f_lw_axi_master_rready
	wire   [3:0] cpu_h2f_lw_axi_master_awlen;                  // cpu:h2f_lw_AWLEN -> mm_interconnect_1:cpu_h2f_lw_axi_master_awlen
	wire  [11:0] cpu_h2f_lw_axi_master_wid;                    // cpu:h2f_lw_WID -> mm_interconnect_1:cpu_h2f_lw_axi_master_wid
	wire   [3:0] cpu_h2f_lw_axi_master_arcache;                // cpu:h2f_lw_ARCACHE -> mm_interconnect_1:cpu_h2f_lw_axi_master_arcache
	wire         cpu_h2f_lw_axi_master_wvalid;                 // cpu:h2f_lw_WVALID -> mm_interconnect_1:cpu_h2f_lw_axi_master_wvalid
	wire  [20:0] cpu_h2f_lw_axi_master_araddr;                 // cpu:h2f_lw_ARADDR -> mm_interconnect_1:cpu_h2f_lw_axi_master_araddr
	wire   [2:0] cpu_h2f_lw_axi_master_arprot;                 // cpu:h2f_lw_ARPROT -> mm_interconnect_1:cpu_h2f_lw_axi_master_arprot
	wire   [2:0] cpu_h2f_lw_axi_master_awprot;                 // cpu:h2f_lw_AWPROT -> mm_interconnect_1:cpu_h2f_lw_axi_master_awprot
	wire  [31:0] cpu_h2f_lw_axi_master_wdata;                  // cpu:h2f_lw_WDATA -> mm_interconnect_1:cpu_h2f_lw_axi_master_wdata
	wire         cpu_h2f_lw_axi_master_arvalid;                // cpu:h2f_lw_ARVALID -> mm_interconnect_1:cpu_h2f_lw_axi_master_arvalid
	wire   [3:0] cpu_h2f_lw_axi_master_awcache;                // cpu:h2f_lw_AWCACHE -> mm_interconnect_1:cpu_h2f_lw_axi_master_awcache
	wire  [11:0] cpu_h2f_lw_axi_master_arid;                   // cpu:h2f_lw_ARID -> mm_interconnect_1:cpu_h2f_lw_axi_master_arid
	wire   [1:0] cpu_h2f_lw_axi_master_arlock;                 // cpu:h2f_lw_ARLOCK -> mm_interconnect_1:cpu_h2f_lw_axi_master_arlock
	wire   [1:0] cpu_h2f_lw_axi_master_awlock;                 // cpu:h2f_lw_AWLOCK -> mm_interconnect_1:cpu_h2f_lw_axi_master_awlock
	wire  [20:0] cpu_h2f_lw_axi_master_awaddr;                 // cpu:h2f_lw_AWADDR -> mm_interconnect_1:cpu_h2f_lw_axi_master_awaddr
	wire   [1:0] cpu_h2f_lw_axi_master_bresp;                  // mm_interconnect_1:cpu_h2f_lw_axi_master_bresp -> cpu:h2f_lw_BRESP
	wire         cpu_h2f_lw_axi_master_arready;                // mm_interconnect_1:cpu_h2f_lw_axi_master_arready -> cpu:h2f_lw_ARREADY
	wire  [31:0] cpu_h2f_lw_axi_master_rdata;                  // mm_interconnect_1:cpu_h2f_lw_axi_master_rdata -> cpu:h2f_lw_RDATA
	wire         cpu_h2f_lw_axi_master_awready;                // mm_interconnect_1:cpu_h2f_lw_axi_master_awready -> cpu:h2f_lw_AWREADY
	wire   [1:0] cpu_h2f_lw_axi_master_arburst;                // cpu:h2f_lw_ARBURST -> mm_interconnect_1:cpu_h2f_lw_axi_master_arburst
	wire   [2:0] cpu_h2f_lw_axi_master_arsize;                 // cpu:h2f_lw_ARSIZE -> mm_interconnect_1:cpu_h2f_lw_axi_master_arsize
	wire         cpu_h2f_lw_axi_master_bready;                 // cpu:h2f_lw_BREADY -> mm_interconnect_1:cpu_h2f_lw_axi_master_bready
	wire         cpu_h2f_lw_axi_master_rlast;                  // mm_interconnect_1:cpu_h2f_lw_axi_master_rlast -> cpu:h2f_lw_RLAST
	wire         cpu_h2f_lw_axi_master_wlast;                  // cpu:h2f_lw_WLAST -> mm_interconnect_1:cpu_h2f_lw_axi_master_wlast
	wire   [1:0] cpu_h2f_lw_axi_master_rresp;                  // mm_interconnect_1:cpu_h2f_lw_axi_master_rresp -> cpu:h2f_lw_RRESP
	wire  [11:0] cpu_h2f_lw_axi_master_awid;                   // cpu:h2f_lw_AWID -> mm_interconnect_1:cpu_h2f_lw_axi_master_awid
	wire  [11:0] cpu_h2f_lw_axi_master_bid;                    // mm_interconnect_1:cpu_h2f_lw_axi_master_bid -> cpu:h2f_lw_BID
	wire         cpu_h2f_lw_axi_master_bvalid;                 // mm_interconnect_1:cpu_h2f_lw_axi_master_bvalid -> cpu:h2f_lw_BVALID
	wire   [2:0] cpu_h2f_lw_axi_master_awsize;                 // cpu:h2f_lw_AWSIZE -> mm_interconnect_1:cpu_h2f_lw_axi_master_awsize
	wire         cpu_h2f_lw_axi_master_awvalid;                // cpu:h2f_lw_AWVALID -> mm_interconnect_1:cpu_h2f_lw_axi_master_awvalid
	wire         cpu_h2f_lw_axi_master_rvalid;                 // mm_interconnect_1:cpu_h2f_lw_axi_master_rvalid -> cpu:h2f_lw_RVALID
	wire         mm_interconnect_1_pio_led_s1_chipselect;      // mm_interconnect_1:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_1_pio_led_s1_readdata;        // pio_led:readdata -> mm_interconnect_1:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_led_s1_address;         // mm_interconnect_1:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_1_pio_led_s1_write;           // mm_interconnect_1:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_1_pio_led_s1_writedata;       // mm_interconnect_1:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_1_pio_display_s1_chipselect;  // mm_interconnect_1:pio_display_s1_chipselect -> pio_display:chipselect
	wire  [31:0] mm_interconnect_1_pio_display_s1_readdata;    // pio_display:readdata -> mm_interconnect_1:pio_display_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_display_s1_address;     // mm_interconnect_1:pio_display_s1_address -> pio_display:address
	wire         mm_interconnect_1_pio_display_s1_write;       // mm_interconnect_1:pio_display_s1_write -> pio_display:write_n
	wire  [31:0] mm_interconnect_1_pio_display_s1_writedata;   // mm_interconnect_1:pio_display_s1_writedata -> pio_display:writedata
	wire         mm_interconnect_1_pio_keys_s1_chipselect;     // mm_interconnect_1:pio_keys_s1_chipselect -> pio_keys:chipselect
	wire  [31:0] mm_interconnect_1_pio_keys_s1_readdata;       // pio_keys:readdata -> mm_interconnect_1:pio_keys_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_keys_s1_address;        // mm_interconnect_1:pio_keys_s1_address -> pio_keys:address
	wire         mm_interconnect_1_pio_keys_s1_write;          // mm_interconnect_1:pio_keys_s1_write -> pio_keys:write_n
	wire  [31:0] mm_interconnect_1_pio_keys_s1_writedata;      // mm_interconnect_1:pio_keys_s1_writedata -> pio_keys:writedata
	wire  [31:0] mm_interconnect_1_pio_fpga2hps_s1_readdata;   // pio_fpga2hps:readdata -> mm_interconnect_1:pio_fpga2hps_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_fpga2hps_s1_address;    // mm_interconnect_1:pio_fpga2hps_s1_address -> pio_fpga2hps:address
	wire         mm_interconnect_1_pio_hps2fpga_s1_chipselect; // mm_interconnect_1:pio_hps2fpga_s1_chipselect -> pio_hps2fpga:chipselect
	wire  [31:0] mm_interconnect_1_pio_hps2fpga_s1_readdata;   // pio_hps2fpga:readdata -> mm_interconnect_1:pio_hps2fpga_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_hps2fpga_s1_address;    // mm_interconnect_1:pio_hps2fpga_s1_address -> pio_hps2fpga:address
	wire         mm_interconnect_1_pio_hps2fpga_s1_write;      // mm_interconnect_1:pio_hps2fpga_s1_write -> pio_hps2fpga:write_n
	wire  [31:0] mm_interconnect_1_pio_hps2fpga_s1_writedata;  // mm_interconnect_1:pio_hps2fpga_s1_writedata -> pio_hps2fpga:writedata
	wire         rst_controller_reset_out_reset;               // rst_controller:reset_out -> [mm_interconnect_0:ram_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:pio_led_reset_reset_bridge_in_reset_reset, pio_display:reset_n, pio_fpga2hps:reset_n, pio_hps2fpga:reset_n, pio_keys:reset_n, pio_led:reset_n, ram:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;           // rst_controller:reset_req -> [ram:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;           // rst_controller_001:reset_out -> [mm_interconnect_0:cpu_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire         cpu_h2f_reset_reset;                          // cpu:h2f_rst_n -> rst_controller_001:reset_in0

	arm_hps_cpu #(
		.F2S_Width (1),
		.S2F_Width (1)
	) cpu (
		.mem_a              (memory_mem_a),                  //            memory.mem_a
		.mem_ba             (memory_mem_ba),                 //                  .mem_ba
		.mem_ck             (memory_mem_ck),                 //                  .mem_ck
		.mem_ck_n           (memory_mem_ck_n),               //                  .mem_ck_n
		.mem_cke            (memory_mem_cke),                //                  .mem_cke
		.mem_cs_n           (memory_mem_cs_n),               //                  .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),              //                  .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),              //                  .mem_cas_n
		.mem_we_n           (memory_mem_we_n),               //                  .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),            //                  .mem_reset_n
		.mem_dq             (memory_mem_dq),                 //                  .mem_dq
		.mem_dqs            (memory_mem_dqs),                //                  .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),              //                  .mem_dqs_n
		.mem_odt            (memory_mem_odt),                //                  .mem_odt
		.mem_dm             (memory_mem_dm),                 //                  .mem_dm
		.oct_rzqin          (memory_oct_rzqin),              //                  .oct_rzqin
		.h2f_rst_n          (cpu_h2f_reset_reset),           //         h2f_reset.reset_n
		.f2h_sdram0_clk     (clk_clk),                       //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR  (),                              //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN   (),                              //                  .arlen
		.f2h_sdram0_ARID    (),                              //                  .arid
		.f2h_sdram0_ARSIZE  (),                              //                  .arsize
		.f2h_sdram0_ARBURST (),                              //                  .arburst
		.f2h_sdram0_ARLOCK  (),                              //                  .arlock
		.f2h_sdram0_ARPROT  (),                              //                  .arprot
		.f2h_sdram0_ARVALID (),                              //                  .arvalid
		.f2h_sdram0_ARCACHE (),                              //                  .arcache
		.f2h_sdram0_AWADDR  (),                              //                  .awaddr
		.f2h_sdram0_AWLEN   (),                              //                  .awlen
		.f2h_sdram0_AWID    (),                              //                  .awid
		.f2h_sdram0_AWSIZE  (),                              //                  .awsize
		.f2h_sdram0_AWBURST (),                              //                  .awburst
		.f2h_sdram0_AWLOCK  (),                              //                  .awlock
		.f2h_sdram0_AWPROT  (),                              //                  .awprot
		.f2h_sdram0_AWVALID (),                              //                  .awvalid
		.f2h_sdram0_AWCACHE (),                              //                  .awcache
		.f2h_sdram0_BRESP   (),                              //                  .bresp
		.f2h_sdram0_BID     (),                              //                  .bid
		.f2h_sdram0_BVALID  (),                              //                  .bvalid
		.f2h_sdram0_BREADY  (),                              //                  .bready
		.f2h_sdram0_ARREADY (),                              //                  .arready
		.f2h_sdram0_AWREADY (),                              //                  .awready
		.f2h_sdram0_RREADY  (),                              //                  .rready
		.f2h_sdram0_RDATA   (),                              //                  .rdata
		.f2h_sdram0_RRESP   (),                              //                  .rresp
		.f2h_sdram0_RLAST   (),                              //                  .rlast
		.f2h_sdram0_RID     (),                              //                  .rid
		.f2h_sdram0_RVALID  (),                              //                  .rvalid
		.f2h_sdram0_WLAST   (),                              //                  .wlast
		.f2h_sdram0_WVALID  (),                              //                  .wvalid
		.f2h_sdram0_WDATA   (),                              //                  .wdata
		.f2h_sdram0_WSTRB   (),                              //                  .wstrb
		.f2h_sdram0_WREADY  (),                              //                  .wready
		.f2h_sdram0_WID     (),                              //                  .wid
		.h2f_axi_clk        (clk_clk),                       //     h2f_axi_clock.clk
		.h2f_AWID           (cpu_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR         (cpu_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN          (cpu_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE         (cpu_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST        (cpu_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK         (cpu_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE        (cpu_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT         (cpu_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID        (cpu_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY        (cpu_h2f_axi_master_awready),    //                  .awready
		.h2f_WID            (cpu_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA          (cpu_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB          (cpu_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST          (cpu_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID         (cpu_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY         (cpu_h2f_axi_master_wready),     //                  .wready
		.h2f_BID            (cpu_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP          (cpu_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID         (cpu_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY         (cpu_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID           (cpu_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR         (cpu_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN          (cpu_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE         (cpu_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST        (cpu_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK         (cpu_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE        (cpu_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT         (cpu_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID        (cpu_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY        (cpu_h2f_axi_master_arready),    //                  .arready
		.h2f_RID            (cpu_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA          (cpu_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP          (cpu_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST          (cpu_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID         (cpu_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY         (cpu_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk        (clk_clk),                       //     f2h_axi_clock.clk
		.f2h_AWID           (),                              //     f2h_axi_slave.awid
		.f2h_AWADDR         (),                              //                  .awaddr
		.f2h_AWLEN          (),                              //                  .awlen
		.f2h_AWSIZE         (),                              //                  .awsize
		.f2h_AWBURST        (),                              //                  .awburst
		.f2h_AWLOCK         (),                              //                  .awlock
		.f2h_AWCACHE        (),                              //                  .awcache
		.f2h_AWPROT         (),                              //                  .awprot
		.f2h_AWVALID        (),                              //                  .awvalid
		.f2h_AWREADY        (),                              //                  .awready
		.f2h_AWUSER         (),                              //                  .awuser
		.f2h_WID            (),                              //                  .wid
		.f2h_WDATA          (),                              //                  .wdata
		.f2h_WSTRB          (),                              //                  .wstrb
		.f2h_WLAST          (),                              //                  .wlast
		.f2h_WVALID         (),                              //                  .wvalid
		.f2h_WREADY         (),                              //                  .wready
		.f2h_BID            (),                              //                  .bid
		.f2h_BRESP          (),                              //                  .bresp
		.f2h_BVALID         (),                              //                  .bvalid
		.f2h_BREADY         (),                              //                  .bready
		.f2h_ARID           (),                              //                  .arid
		.f2h_ARADDR         (),                              //                  .araddr
		.f2h_ARLEN          (),                              //                  .arlen
		.f2h_ARSIZE         (),                              //                  .arsize
		.f2h_ARBURST        (),                              //                  .arburst
		.f2h_ARLOCK         (),                              //                  .arlock
		.f2h_ARCACHE        (),                              //                  .arcache
		.f2h_ARPROT         (),                              //                  .arprot
		.f2h_ARVALID        (),                              //                  .arvalid
		.f2h_ARREADY        (),                              //                  .arready
		.f2h_ARUSER         (),                              //                  .aruser
		.f2h_RID            (),                              //                  .rid
		.f2h_RDATA          (),                              //                  .rdata
		.f2h_RRESP          (),                              //                  .rresp
		.f2h_RLAST          (),                              //                  .rlast
		.f2h_RVALID         (),                              //                  .rvalid
		.f2h_RREADY         (),                              //                  .rready
		.h2f_lw_axi_clk     (clk_clk),                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID        (cpu_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR      (cpu_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN       (cpu_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE      (cpu_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST     (cpu_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK      (cpu_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE     (cpu_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT      (cpu_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID     (cpu_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY     (cpu_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID         (cpu_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA       (cpu_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB       (cpu_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST       (cpu_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID      (cpu_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY      (cpu_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID         (cpu_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP       (cpu_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID      (cpu_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY      (cpu_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID        (cpu_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR      (cpu_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN       (cpu_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE      (cpu_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST     (cpu_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK      (cpu_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE     (cpu_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT      (cpu_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID     (cpu_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY     (cpu_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID         (cpu_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA       (cpu_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP       (cpu_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST       (cpu_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID      (cpu_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY      (cpu_h2f_lw_axi_master_rready)   //                  .rready
	);

	arm_hps_pio_display pio_display (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_pio_display_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_display_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_display_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_display_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_display_s1_readdata),   //                    .readdata
		.out_port   (pio_display_export)                           // external_connection.export
	);

	arm_hps_pio_fpga2hps pio_fpga2hps (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_pio_fpga2hps_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_pio_fpga2hps_s1_readdata), //                    .readdata
		.in_port  (pio_fpga2hps_export)                         // external_connection.export
	);

	arm_hps_pio_hps2fpga pio_hps2fpga (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_pio_hps2fpga_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_hps2fpga_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_hps2fpga_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_hps2fpga_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_hps2fpga_s1_readdata),   //                    .readdata
		.out_port   (pio_hps2fpga_export)                           // external_connection.export
	);

	arm_hps_pio_keys pio_keys (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_1_pio_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_keys_s1_readdata),   //                    .readdata
		.in_port    (pio_keys_export)                           // external_connection.export
	);

	arm_hps_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	arm_hps_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	arm_hps_mm_interconnect_0 mm_interconnect_0 (
		.cpu_h2f_axi_master_awid                                        (cpu_h2f_axi_master_awid),             //                                       cpu_h2f_axi_master.awid
		.cpu_h2f_axi_master_awaddr                                      (cpu_h2f_axi_master_awaddr),           //                                                         .awaddr
		.cpu_h2f_axi_master_awlen                                       (cpu_h2f_axi_master_awlen),            //                                                         .awlen
		.cpu_h2f_axi_master_awsize                                      (cpu_h2f_axi_master_awsize),           //                                                         .awsize
		.cpu_h2f_axi_master_awburst                                     (cpu_h2f_axi_master_awburst),          //                                                         .awburst
		.cpu_h2f_axi_master_awlock                                      (cpu_h2f_axi_master_awlock),           //                                                         .awlock
		.cpu_h2f_axi_master_awcache                                     (cpu_h2f_axi_master_awcache),          //                                                         .awcache
		.cpu_h2f_axi_master_awprot                                      (cpu_h2f_axi_master_awprot),           //                                                         .awprot
		.cpu_h2f_axi_master_awvalid                                     (cpu_h2f_axi_master_awvalid),          //                                                         .awvalid
		.cpu_h2f_axi_master_awready                                     (cpu_h2f_axi_master_awready),          //                                                         .awready
		.cpu_h2f_axi_master_wid                                         (cpu_h2f_axi_master_wid),              //                                                         .wid
		.cpu_h2f_axi_master_wdata                                       (cpu_h2f_axi_master_wdata),            //                                                         .wdata
		.cpu_h2f_axi_master_wstrb                                       (cpu_h2f_axi_master_wstrb),            //                                                         .wstrb
		.cpu_h2f_axi_master_wlast                                       (cpu_h2f_axi_master_wlast),            //                                                         .wlast
		.cpu_h2f_axi_master_wvalid                                      (cpu_h2f_axi_master_wvalid),           //                                                         .wvalid
		.cpu_h2f_axi_master_wready                                      (cpu_h2f_axi_master_wready),           //                                                         .wready
		.cpu_h2f_axi_master_bid                                         (cpu_h2f_axi_master_bid),              //                                                         .bid
		.cpu_h2f_axi_master_bresp                                       (cpu_h2f_axi_master_bresp),            //                                                         .bresp
		.cpu_h2f_axi_master_bvalid                                      (cpu_h2f_axi_master_bvalid),           //                                                         .bvalid
		.cpu_h2f_axi_master_bready                                      (cpu_h2f_axi_master_bready),           //                                                         .bready
		.cpu_h2f_axi_master_arid                                        (cpu_h2f_axi_master_arid),             //                                                         .arid
		.cpu_h2f_axi_master_araddr                                      (cpu_h2f_axi_master_araddr),           //                                                         .araddr
		.cpu_h2f_axi_master_arlen                                       (cpu_h2f_axi_master_arlen),            //                                                         .arlen
		.cpu_h2f_axi_master_arsize                                      (cpu_h2f_axi_master_arsize),           //                                                         .arsize
		.cpu_h2f_axi_master_arburst                                     (cpu_h2f_axi_master_arburst),          //                                                         .arburst
		.cpu_h2f_axi_master_arlock                                      (cpu_h2f_axi_master_arlock),           //                                                         .arlock
		.cpu_h2f_axi_master_arcache                                     (cpu_h2f_axi_master_arcache),          //                                                         .arcache
		.cpu_h2f_axi_master_arprot                                      (cpu_h2f_axi_master_arprot),           //                                                         .arprot
		.cpu_h2f_axi_master_arvalid                                     (cpu_h2f_axi_master_arvalid),          //                                                         .arvalid
		.cpu_h2f_axi_master_arready                                     (cpu_h2f_axi_master_arready),          //                                                         .arready
		.cpu_h2f_axi_master_rid                                         (cpu_h2f_axi_master_rid),              //                                                         .rid
		.cpu_h2f_axi_master_rdata                                       (cpu_h2f_axi_master_rdata),            //                                                         .rdata
		.cpu_h2f_axi_master_rresp                                       (cpu_h2f_axi_master_rresp),            //                                                         .rresp
		.cpu_h2f_axi_master_rlast                                       (cpu_h2f_axi_master_rlast),            //                                                         .rlast
		.cpu_h2f_axi_master_rvalid                                      (cpu_h2f_axi_master_rvalid),           //                                                         .rvalid
		.cpu_h2f_axi_master_rready                                      (cpu_h2f_axi_master_rready),           //                                                         .rready
		.clk_50mhz_clk_clk                                              (clk_clk),                             //                                            clk_50mhz_clk.clk
		.cpu_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),  // cpu_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.ram_reset1_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),      //                         ram_reset1_reset_bridge_in_reset.reset
		.ram_s1_address                                                 (mm_interconnect_0_ram_s1_address),    //                                                   ram_s1.address
		.ram_s1_write                                                   (mm_interconnect_0_ram_s1_write),      //                                                         .write
		.ram_s1_readdata                                                (mm_interconnect_0_ram_s1_readdata),   //                                                         .readdata
		.ram_s1_writedata                                               (mm_interconnect_0_ram_s1_writedata),  //                                                         .writedata
		.ram_s1_byteenable                                              (mm_interconnect_0_ram_s1_byteenable), //                                                         .byteenable
		.ram_s1_chipselect                                              (mm_interconnect_0_ram_s1_chipselect), //                                                         .chipselect
		.ram_s1_clken                                                   (mm_interconnect_0_ram_s1_clken)       //                                                         .clken
	);

	arm_hps_mm_interconnect_1 mm_interconnect_1 (
		.cpu_h2f_lw_axi_master_awid                                        (cpu_h2f_lw_axi_master_awid),                   //                                       cpu_h2f_lw_axi_master.awid
		.cpu_h2f_lw_axi_master_awaddr                                      (cpu_h2f_lw_axi_master_awaddr),                 //                                                            .awaddr
		.cpu_h2f_lw_axi_master_awlen                                       (cpu_h2f_lw_axi_master_awlen),                  //                                                            .awlen
		.cpu_h2f_lw_axi_master_awsize                                      (cpu_h2f_lw_axi_master_awsize),                 //                                                            .awsize
		.cpu_h2f_lw_axi_master_awburst                                     (cpu_h2f_lw_axi_master_awburst),                //                                                            .awburst
		.cpu_h2f_lw_axi_master_awlock                                      (cpu_h2f_lw_axi_master_awlock),                 //                                                            .awlock
		.cpu_h2f_lw_axi_master_awcache                                     (cpu_h2f_lw_axi_master_awcache),                //                                                            .awcache
		.cpu_h2f_lw_axi_master_awprot                                      (cpu_h2f_lw_axi_master_awprot),                 //                                                            .awprot
		.cpu_h2f_lw_axi_master_awvalid                                     (cpu_h2f_lw_axi_master_awvalid),                //                                                            .awvalid
		.cpu_h2f_lw_axi_master_awready                                     (cpu_h2f_lw_axi_master_awready),                //                                                            .awready
		.cpu_h2f_lw_axi_master_wid                                         (cpu_h2f_lw_axi_master_wid),                    //                                                            .wid
		.cpu_h2f_lw_axi_master_wdata                                       (cpu_h2f_lw_axi_master_wdata),                  //                                                            .wdata
		.cpu_h2f_lw_axi_master_wstrb                                       (cpu_h2f_lw_axi_master_wstrb),                  //                                                            .wstrb
		.cpu_h2f_lw_axi_master_wlast                                       (cpu_h2f_lw_axi_master_wlast),                  //                                                            .wlast
		.cpu_h2f_lw_axi_master_wvalid                                      (cpu_h2f_lw_axi_master_wvalid),                 //                                                            .wvalid
		.cpu_h2f_lw_axi_master_wready                                      (cpu_h2f_lw_axi_master_wready),                 //                                                            .wready
		.cpu_h2f_lw_axi_master_bid                                         (cpu_h2f_lw_axi_master_bid),                    //                                                            .bid
		.cpu_h2f_lw_axi_master_bresp                                       (cpu_h2f_lw_axi_master_bresp),                  //                                                            .bresp
		.cpu_h2f_lw_axi_master_bvalid                                      (cpu_h2f_lw_axi_master_bvalid),                 //                                                            .bvalid
		.cpu_h2f_lw_axi_master_bready                                      (cpu_h2f_lw_axi_master_bready),                 //                                                            .bready
		.cpu_h2f_lw_axi_master_arid                                        (cpu_h2f_lw_axi_master_arid),                   //                                                            .arid
		.cpu_h2f_lw_axi_master_araddr                                      (cpu_h2f_lw_axi_master_araddr),                 //                                                            .araddr
		.cpu_h2f_lw_axi_master_arlen                                       (cpu_h2f_lw_axi_master_arlen),                  //                                                            .arlen
		.cpu_h2f_lw_axi_master_arsize                                      (cpu_h2f_lw_axi_master_arsize),                 //                                                            .arsize
		.cpu_h2f_lw_axi_master_arburst                                     (cpu_h2f_lw_axi_master_arburst),                //                                                            .arburst
		.cpu_h2f_lw_axi_master_arlock                                      (cpu_h2f_lw_axi_master_arlock),                 //                                                            .arlock
		.cpu_h2f_lw_axi_master_arcache                                     (cpu_h2f_lw_axi_master_arcache),                //                                                            .arcache
		.cpu_h2f_lw_axi_master_arprot                                      (cpu_h2f_lw_axi_master_arprot),                 //                                                            .arprot
		.cpu_h2f_lw_axi_master_arvalid                                     (cpu_h2f_lw_axi_master_arvalid),                //                                                            .arvalid
		.cpu_h2f_lw_axi_master_arready                                     (cpu_h2f_lw_axi_master_arready),                //                                                            .arready
		.cpu_h2f_lw_axi_master_rid                                         (cpu_h2f_lw_axi_master_rid),                    //                                                            .rid
		.cpu_h2f_lw_axi_master_rdata                                       (cpu_h2f_lw_axi_master_rdata),                  //                                                            .rdata
		.cpu_h2f_lw_axi_master_rresp                                       (cpu_h2f_lw_axi_master_rresp),                  //                                                            .rresp
		.cpu_h2f_lw_axi_master_rlast                                       (cpu_h2f_lw_axi_master_rlast),                  //                                                            .rlast
		.cpu_h2f_lw_axi_master_rvalid                                      (cpu_h2f_lw_axi_master_rvalid),                 //                                                            .rvalid
		.cpu_h2f_lw_axi_master_rready                                      (cpu_h2f_lw_axi_master_rready),                 //                                                            .rready
		.clk_50mhz_clk_clk                                                 (clk_clk),                                      //                                               clk_50mhz_clk.clk
		.cpu_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),           // cpu_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pio_led_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),               //                         pio_led_reset_reset_bridge_in_reset.reset
		.pio_display_s1_address                                            (mm_interconnect_1_pio_display_s1_address),     //                                              pio_display_s1.address
		.pio_display_s1_write                                              (mm_interconnect_1_pio_display_s1_write),       //                                                            .write
		.pio_display_s1_readdata                                           (mm_interconnect_1_pio_display_s1_readdata),    //                                                            .readdata
		.pio_display_s1_writedata                                          (mm_interconnect_1_pio_display_s1_writedata),   //                                                            .writedata
		.pio_display_s1_chipselect                                         (mm_interconnect_1_pio_display_s1_chipselect),  //                                                            .chipselect
		.pio_fpga2hps_s1_address                                           (mm_interconnect_1_pio_fpga2hps_s1_address),    //                                             pio_fpga2hps_s1.address
		.pio_fpga2hps_s1_readdata                                          (mm_interconnect_1_pio_fpga2hps_s1_readdata),   //                                                            .readdata
		.pio_hps2fpga_s1_address                                           (mm_interconnect_1_pio_hps2fpga_s1_address),    //                                             pio_hps2fpga_s1.address
		.pio_hps2fpga_s1_write                                             (mm_interconnect_1_pio_hps2fpga_s1_write),      //                                                            .write
		.pio_hps2fpga_s1_readdata                                          (mm_interconnect_1_pio_hps2fpga_s1_readdata),   //                                                            .readdata
		.pio_hps2fpga_s1_writedata                                         (mm_interconnect_1_pio_hps2fpga_s1_writedata),  //                                                            .writedata
		.pio_hps2fpga_s1_chipselect                                        (mm_interconnect_1_pio_hps2fpga_s1_chipselect), //                                                            .chipselect
		.pio_keys_s1_address                                               (mm_interconnect_1_pio_keys_s1_address),        //                                                 pio_keys_s1.address
		.pio_keys_s1_write                                                 (mm_interconnect_1_pio_keys_s1_write),          //                                                            .write
		.pio_keys_s1_readdata                                              (mm_interconnect_1_pio_keys_s1_readdata),       //                                                            .readdata
		.pio_keys_s1_writedata                                             (mm_interconnect_1_pio_keys_s1_writedata),      //                                                            .writedata
		.pio_keys_s1_chipselect                                            (mm_interconnect_1_pio_keys_s1_chipselect),     //                                                            .chipselect
		.pio_led_s1_address                                                (mm_interconnect_1_pio_led_s1_address),         //                                                  pio_led_s1.address
		.pio_led_s1_write                                                  (mm_interconnect_1_pio_led_s1_write),           //                                                            .write
		.pio_led_s1_readdata                                               (mm_interconnect_1_pio_led_s1_readdata),        //                                                            .readdata
		.pio_led_s1_writedata                                              (mm_interconnect_1_pio_led_s1_writedata),       //                                                            .writedata
		.pio_led_s1_chipselect                                             (mm_interconnect_1_pio_led_s1_chipselect)       //                                                            .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~cpu_h2f_reset_reset),               // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
